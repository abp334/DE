<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>4.55849,-0.136664,107.833,-51.1835</PageViewport>
<gate>
<ID>2</ID>
<type>AA_MUX_2x1</type>
<position>31.5,-15</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>4 </output>
<input>
<ID>SEL_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>23.5,-14</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>23.5,-17</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>28,-10.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>36.5,-15</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>26.5,-24</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>20.5,-34.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>19,-28</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>48.5,-22.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_INVERTER</type>
<position>33,-27.5</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>36.5,-32</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_OR2</type>
<position>55.5,-28</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>GA_LED</type>
<position>60.5,-28</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>46,-14</position>
<gparam>LABEL_TEXT 2x1 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>36.5,-37.5</position>
<gparam>LABEL_TEXT Using AOI logic</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-14,29.5,-14</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>29.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>29.5,-14,29.5,-14</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-14 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-17,27.5,-16</points>
<intersection>-17 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-16,29.5,-16</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-17,27.5,-17</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-12.5,31.5,-10.5</points>
<connection>
<GID>2</GID>
<name>SEL_0</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-10.5,31.5,-10.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-15,35.5,-15</points>
<connection>
<GID>10</GID>
<name>N_in0</name></connection>
<connection>
<GID>2</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21,-27.5,30,-27.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>21 4</intersection>
<intersection>25 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>21,-28,21,-27.5</points>
<intersection>-28 7</intersection>
<intersection>-27.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>25,-31,25,-27.5</points>
<intersection>-31 6</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>25,-31,33.5,-31</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>25 5</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>21,-28,21,-28</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>21 4</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-27.5,36,-23.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-23.5,45.5,-23.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-24,32.5,-21.5</points>
<intersection>-24 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-21.5,45.5,-21.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-24,32.5,-24</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-34.5,32,-33</points>
<intersection>-34.5 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-33,33.5,-33</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-34.5,32,-34.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-27,52,-22.5</points>
<intersection>-27 1</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-27,52.5,-27</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-22.5,52,-22.5</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-32,46,-29</points>
<intersection>-32 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-29,52.5,-29</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39.5,-32,46,-32</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-28,59.5,-28</points>
<connection>
<GID>26</GID>
<name>N_in0</name></connection>
<connection>
<GID>24</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>21.6705,6.8864,113.471,-38.4886</PageViewport>
<gate>
<ID>32</ID>
<type>AE_MUX_4x1</type>
<position>47,-16</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>13 </input>
<input>
<ID>IN_3</ID>12 </input>
<output>
<ID>OUT</ID>18 </output>
<input>
<ID>SEL_0</ID>17 </input>
<input>
<ID>SEL_1</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>35.5,-13</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>35.5,-15.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>35.5,-18</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>35.5,-20.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>42,-8</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>42,-5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>46</ID>
<type>GA_LED</type>
<position>52,-16</position>
<input>
<ID>N_in0</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>48,-23.5</position>
<gparam>LABEL_TEXT 4x1 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-13,44,-13</points>
<connection>
<GID>32</GID>
<name>IN_3</name></connection>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-15.5,40.5,-15</points>
<intersection>-15.5 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-15,44,-15</points>
<connection>
<GID>32</GID>
<name>IN_2</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-15.5,40.5,-15.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-18,40.5,-17</points>
<intersection>-18 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-17,44,-17</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-18,40.5,-18</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-20.5,40.5,-19</points>
<intersection>-20.5 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-19,44,-19</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-20.5,40.5,-20.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-11,47,-8</points>
<connection>
<GID>32</GID>
<name>SEL_1</name></connection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-8,47,-8</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-11,48,-5</points>
<connection>
<GID>32</GID>
<name>SEL_0</name></connection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-5,48,-5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-16,51,-16</points>
<connection>
<GID>46</GID>
<name>N_in0</name></connection>
<connection>
<GID>32</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>7.38751,-4.68125,99.1875,-50.0563</PageViewport>
<gate>
<ID>48</ID>
<type>BA_DECODER_2x4</type>
<position>40.5,-21.5</position>
<input>
<ID>ENABLE</ID>19 </input>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT_0</ID>25 </output>
<output>
<ID>OUT_1</ID>24 </output>
<output>
<ID>OUT_2</ID>23 </output>
<output>
<ID>OUT_3</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>32,-20</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_TOGGLE</type>
<position>32,-22.5</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_TOGGLE</type>
<position>32,-25</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>56</ID>
<type>GA_LED</type>
<position>47,-19.5</position>
<input>
<ID>N_in0</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>GA_LED</type>
<position>54.5,-21</position>
<input>
<ID>N_in0</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>GA_LED</type>
<position>53,-23.5</position>
<input>
<ID>N_in0</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>GA_LED</type>
<position>47,-28</position>
<input>
<ID>N_in0</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>38.5,-31</position>
<gparam>LABEL_TEXT 2x4 Decoder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-20,37.5,-20</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>37.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37.5,-20,37.5,-20</points>
<connection>
<GID>48</GID>
<name>ENABLE</name></connection>
<intersection>-20 1</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-22.5,35.5,-22</points>
<intersection>-22.5 2</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-22,37.5,-22</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-22.5,35.5,-22.5</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-25,35.5,-23</points>
<intersection>-25 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-23,37.5,-23</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-25,35.5,-25</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-20,44.5,-19.5</points>
<intersection>-20 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-19.5,46,-19.5</points>
<connection>
<GID>56</GID>
<name>N_in0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-20,44.5,-20</points>
<connection>
<GID>48</GID>
<name>OUT_3</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43.5,-21,53.5,-21</points>
<connection>
<GID>48</GID>
<name>OUT_2</name></connection>
<connection>
<GID>58</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-23.5,44.5,-22</points>
<intersection>-23.5 1</intersection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-23.5,52,-23.5</points>
<connection>
<GID>60</GID>
<name>N_in0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-22,44.5,-22</points>
<connection>
<GID>48</GID>
<name>OUT_1</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-28,43.5,-23</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-28,46,-28</points>
<connection>
<GID>64</GID>
<name>N_in0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport>
<gate>
<ID>70</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>42,-22</position>
<output>
<ID>A_equal_B</ID>41 </output>
<output>
<ID>A_greater_B</ID>40 </output>
<output>
<ID>A_less_B</ID>42 </output>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>30 </input>
<input>
<ID>IN_2</ID>28 </input>
<input>
<ID>IN_3</ID>27 </input>
<input>
<ID>IN_B_0</ID>32 </input>
<input>
<ID>IN_B_1</ID>33 </input>
<input>
<ID>IN_B_2</ID>34 </input>
<input>
<ID>IN_B_3</ID>35 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>31,-14.5</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_TOGGLE</type>
<position>31,-11.5</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_TOGGLE</type>
<position>31,-8.5</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_TOGGLE</type>
<position>31,-5.5</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_TOGGLE</type>
<position>53,-15</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_TOGGLE</type>
<position>53,-12</position>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_TOGGLE</type>
<position>53,-9</position>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_TOGGLE</type>
<position>53,-6</position>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>94</ID>
<type>GA_LED</type>
<position>29.5,-20</position>
<input>
<ID>N_in1</ID>40 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>GA_LED</type>
<position>29.5,-22.5</position>
<input>
<ID>N_in1</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>GA_LED</type>
<position>29.5,-25.5</position>
<input>
<ID>N_in1</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>AA_LABEL</type>
<position>43.5,-28</position>
<gparam>LABEL_TEXT Comparator</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-18,37,-14.5</points>
<connection>
<GID>70</GID>
<name>IN_3</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-14.5,37,-14.5</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-18,38,-11.5</points>
<connection>
<GID>70</GID>
<name>IN_2</name></connection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-11.5,38,-11.5</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-18,39,-8.5</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-8.5,39,-8.5</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-18,40,-5.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-5.5,40,-5.5</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-18,47,-15</points>
<connection>
<GID>70</GID>
<name>IN_B_0</name></connection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>47,-15,51,-15</points>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-18,46,-12</points>
<connection>
<GID>70</GID>
<name>IN_B_1</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-12,51,-12</points>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-18,45,-9</points>
<connection>
<GID>70</GID>
<name>IN_B_2</name></connection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-9,51,-9</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-18,44,-6</points>
<connection>
<GID>70</GID>
<name>IN_B_3</name></connection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-6,51,-6</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-20,34,-20</points>
<connection>
<GID>70</GID>
<name>A_greater_B</name></connection>
<connection>
<GID>94</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-22.5,32,-22</points>
<intersection>-22.5 2</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-22,34,-22</points>
<connection>
<GID>70</GID>
<name>A_equal_B</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-22.5,32,-22.5</points>
<connection>
<GID>96</GID>
<name>N_in1</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-25.5,32,-24</points>
<intersection>-25.5 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-24,34,-24</points>
<connection>
<GID>70</GID>
<name>A_less_B</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-25.5,32,-25.5</points>
<connection>
<GID>98</GID>
<name>N_in1</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>20.1,0.799999,142.5,-59.7</PageViewport>
<gate>
<ID>102</ID>
<type>AI_XOR2</type>
<position>48.5,-16</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>AI_XOR2</type>
<position>49,-24.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>108</ID>
<type>AI_XOR2</type>
<position>49.5,-35</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_TOGGLE</type>
<position>34.5,-12</position>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_TOGGLE</type>
<position>34.5,-18</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>114</ID>
<type>AA_TOGGLE</type>
<position>34,-25</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>116</ID>
<type>AA_TOGGLE</type>
<position>33.5,-36</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>118</ID>
<type>GA_LED</type>
<position>56,-11.5</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>GA_LED</type>
<position>54.5,-16</position>
<input>
<ID>N_in0</ID>47 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>GA_LED</type>
<position>54.5,-24.5</position>
<input>
<ID>N_in0</ID>48 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>GA_LED</type>
<position>54.5,-35</position>
<input>
<ID>N_in0</ID>49 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>45.5,-41</position>
<gparam>LABEL_TEXT 4-bit Binary to Gray converter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>AI_XOR2</type>
<position>92,-13</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>51 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>130</ID>
<type>AI_XOR2</type>
<position>101,-23.5</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>52 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>132</ID>
<type>AI_XOR2</type>
<position>113.5,-33.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>53 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>AA_TOGGLE</type>
<position>80,-10</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>136</ID>
<type>AA_TOGGLE</type>
<position>80,-14</position>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>138</ID>
<type>AA_TOGGLE</type>
<position>79.5,-21.5</position>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>140</ID>
<type>AA_TOGGLE</type>
<position>79.5,-30</position>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>142</ID>
<type>GA_LED</type>
<position>100.5,-10</position>
<input>
<ID>N_in0</ID>50 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>144</ID>
<type>GA_LED</type>
<position>101,-13</position>
<input>
<ID>N_in0</ID>54 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>146</ID>
<type>GA_LED</type>
<position>113,-23.5</position>
<input>
<ID>N_in0</ID>55 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>GA_LED</type>
<position>118.5,-33.5</position>
<input>
<ID>N_in0</ID>56 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>AA_LABEL</type>
<position>101,-41</position>
<gparam>LABEL_TEXT 4-bit Gray to Binary converter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36.5,-12,55,-12</points>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection>
<intersection>45.5 4</intersection>
<intersection>55 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>55,-12,55,-11.5</points>
<connection>
<GID>118</GID>
<name>N_in0</name></connection>
<intersection>-12 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>45.5,-15,45.5,-12</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>-12 1</intersection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36.5,-17,45.5,-17</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>36.5 5</intersection>
<intersection>42.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>42.5,-23.5,42.5,-17</points>
<intersection>-23.5 4</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>42.5,-23.5,46,-23.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>42.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>36.5,-18,36.5,-17</points>
<connection>
<GID>112</GID>
<name>OUT_0</name></connection>
<intersection>-17 1</intersection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-25.5,46,-25.5</points>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>36 3</intersection>
<intersection>41 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36,-25.5,36,-25</points>
<connection>
<GID>114</GID>
<name>OUT_0</name></connection>
<intersection>-25.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>41,-34,41,-25.5</points>
<intersection>-34 5</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>41,-34,46.5,-34</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>41 4</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-36,46.5,-36</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<connection>
<GID>116</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51.5,-16,53.5,-16</points>
<connection>
<GID>120</GID>
<name>N_in0</name></connection>
<connection>
<GID>102</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52,-24.5,53.5,-24.5</points>
<connection>
<GID>122</GID>
<name>N_in0</name></connection>
<connection>
<GID>106</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52.5,-35,53.5,-35</points>
<connection>
<GID>124</GID>
<name>N_in0</name></connection>
<connection>
<GID>108</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82,-10,99.5,-10</points>
<connection>
<GID>142</GID>
<name>N_in0</name></connection>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection>
<intersection>89 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>89,-12,89,-10</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>-10 1</intersection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82,-14,89,-14</points>
<connection>
<GID>128</GID>
<name>IN_1</name></connection>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81.5,-24.5,98,-24.5</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>81.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>81.5,-24.5,81.5,-21.5</points>
<connection>
<GID>138</GID>
<name>OUT_0</name></connection>
<intersection>-24.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81.5,-34.5,110.5,-34.5</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<intersection>81.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>81.5,-34.5,81.5,-30</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<intersection>-34.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>95,-13,100,-13</points>
<connection>
<GID>128</GID>
<name>OUT</name></connection>
<connection>
<GID>144</GID>
<name>N_in0</name></connection>
<intersection>97 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>97,-22.5,97,-13</points>
<intersection>-22.5 4</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>97,-22.5,98,-22.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>97 3</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104,-23.5,112,-23.5</points>
<connection>
<GID>130</GID>
<name>OUT</name></connection>
<connection>
<GID>146</GID>
<name>N_in0</name></connection>
<intersection>108 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>108,-32.5,108,-23.5</points>
<intersection>-32.5 7</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>108,-32.5,110.5,-32.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>108 6</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116.5,-33.5,117.5,-33.5</points>
<connection>
<GID>148</GID>
<name>N_in0</name></connection>
<connection>
<GID>132</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport>
<gate>
<ID>212</ID>
<type>AA_LABEL</type>
<position>24,-27</position>
<gparam>LABEL_TEXT D-FLIPFLOP</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>AE_DFF_LOW</type>
<position>50.5,-11</position>
<input>
<ID>IN_0</ID>64 </input>
<output>
<ID>OUTINV_0</ID>69 </output>
<output>
<ID>OUT_0</ID>68 </output>
<input>
<ID>clock</ID>67 </input>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>164</ID>
<type>DA_FROM</type>
<position>42.5,-9</position>
<input>
<ID>IN_0</ID>64 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>166</ID>
<type>DE_TO</type>
<position>28,-13</position>
<input>
<ID>IN_0</ID>65 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>168</ID>
<type>AA_TOGGLE</type>
<position>23,-16</position>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>170</ID>
<type>BB_CLOCK</type>
<position>46,-30</position>
<output>
<ID>CLK</ID>66 </output>
<gparam>angle 0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>172</ID>
<type>DA_FROM</type>
<position>42.5,-12</position>
<input>
<ID>IN_0</ID>67 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>174</ID>
<type>DE_TO</type>
<position>55.5,-30</position>
<input>
<ID>IN_0</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>176</ID>
<type>GA_LED</type>
<position>56,-9</position>
<input>
<ID>N_in0</ID>68 </input>
<input>
<ID>N_in1</ID>70 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>GA_LED</type>
<position>56,-12</position>
<input>
<ID>N_in0</ID>69 </input>
<input>
<ID>N_in1</ID>71 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>180</ID>
<type>DE_TO</type>
<position>62.5,-9</position>
<input>
<ID>IN_0</ID>70 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q</lparam></gate>
<gate>
<ID>182</ID>
<type>DE_TO</type>
<position>60.5,-12</position>
<input>
<ID>IN_0</ID>71 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q'</lparam></gate>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44.5,-9,47.5,-9</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>47.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>47.5,-9,47.5,-9</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>-9 1</intersection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-14,23,-13</points>
<connection>
<GID>168</GID>
<name>OUT_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-13,26,-13</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-30,53.5,-30</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>50 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>50,-30,50,-30</points>
<connection>
<GID>170</GID>
<name>CLK</name></connection>
<intersection>-30 1</intersection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44.5,-12,47.5,-12</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>47.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>47.5,-12,47.5,-12</points>
<connection>
<GID>152</GID>
<name>clock</name></connection>
<intersection>-12 1</intersection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-9,55,-9</points>
<connection>
<GID>176</GID>
<name>N_in0</name></connection>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-12,55,-12</points>
<connection>
<GID>152</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>178</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-9,60.5,-9</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>57 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>57,-9,57,-9</points>
<connection>
<GID>176</GID>
<name>N_in1</name></connection>
<intersection>-9 1</intersection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-12,58.5,-12</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>57 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>57,-12,57,-12</points>
<connection>
<GID>178</GID>
<name>N_in1</name></connection>
<intersection>-12 1</intersection></vsegment></shape></wire></page 5>
<page 6>
<PageViewport>4.01875,8.99375,126.419,-51.5063</PageViewport>
<gate>
<ID>194</ID>
<type>GA_LED</type>
<position>56,-18</position>
<input>
<ID>N_in0</ID>76 </input>
<input>
<ID>N_in1</ID>81 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>196</ID>
<type>DE_TO</type>
<position>23.5,-20.5</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID J</lparam></gate>
<gate>
<ID>198</ID>
<type>DE_TO</type>
<position>24,-28.5</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID K</lparam></gate>
<gate>
<ID>200</ID>
<type>DE_TO</type>
<position>25,-37</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK1</lparam></gate>
<gate>
<ID>202</ID>
<type>AA_TOGGLE</type>
<position>17.5,-20.5</position>
<output>
<ID>OUT_0</ID>77 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>204</ID>
<type>AA_TOGGLE</type>
<position>17.5,-28.5</position>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>206</ID>
<type>BB_CLOCK</type>
<position>16.5,-37</position>
<output>
<ID>CLK</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>208</ID>
<type>DE_TO</type>
<position>68,-14</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q1</lparam></gate>
<gate>
<ID>210</ID>
<type>DE_TO</type>
<position>67.5,-18</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q'1</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_LABEL</type>
<position>54.5,-28</position>
<gparam>LABEL_TEXT JK-FLIPFLOP</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>184</ID>
<type>BE_JKFF_LOW</type>
<position>52,-16</position>
<input>
<ID>J</ID>72 </input>
<input>
<ID>K</ID>74 </input>
<output>
<ID>Q</ID>75 </output>
<input>
<ID>clock</ID>73 </input>
<output>
<ID>nQ</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>186</ID>
<type>DA_FROM</type>
<position>38,-14</position>
<input>
<ID>IN_0</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID J</lparam></gate>
<gate>
<ID>188</ID>
<type>DA_FROM</type>
<position>44,-16</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK1</lparam></gate>
<gate>
<ID>190</ID>
<type>DA_FROM</type>
<position>38.5,-18</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID K</lparam></gate>
<gate>
<ID>192</ID>
<type>GA_LED</type>
<position>56,-14</position>
<input>
<ID>N_in0</ID>75 </input>
<input>
<ID>N_in1</ID>80 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-14,49,-14</points>
<connection>
<GID>184</GID>
<name>J</name></connection>
<connection>
<GID>186</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46,-16,49,-16</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>49 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>49,-16,49,-16</points>
<connection>
<GID>184</GID>
<name>clock</name></connection>
<intersection>-16 1</intersection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-18,49,-18</points>
<connection>
<GID>184</GID>
<name>K</name></connection>
<connection>
<GID>190</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-14,55,-14</points>
<connection>
<GID>192</GID>
<name>N_in0</name></connection>
<connection>
<GID>184</GID>
<name>Q</name></connection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-18,55,-18</points>
<connection>
<GID>194</GID>
<name>N_in0</name></connection>
<connection>
<GID>184</GID>
<name>nQ</name></connection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-20.5,21.5,-20.5</points>
<connection>
<GID>202</GID>
<name>OUT_0</name></connection>
<intersection>21.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>21.5,-20.5,21.5,-20.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>-20.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-28.5,22,-28.5</points>
<connection>
<GID>204</GID>
<name>OUT_0</name></connection>
<connection>
<GID>198</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-37,23,-37</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>20.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>20.5,-37,20.5,-37</points>
<connection>
<GID>206</GID>
<name>CLK</name></connection>
<intersection>-37 1</intersection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-14,66,-14</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>57 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57,-14,57,-14</points>
<connection>
<GID>192</GID>
<name>N_in1</name></connection>
<intersection>-14 1</intersection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-18,65.5,-18</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<intersection>57 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>57,-18,57,-18</points>
<connection>
<GID>194</GID>
<name>N_in1</name></connection>
<intersection>-18 1</intersection></vsegment></shape></wire></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>