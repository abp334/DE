<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>4.55849,-0.136664,107.833,-51.1835</PageViewport>
<gate>
<ID>2</ID>
<type>AA_MUX_2x1</type>
<position>31.5,-15</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>4 </output>
<input>
<ID>SEL_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>23.5,-14</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>23.5,-17</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>28,-10.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>36.5,-15</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>26.5,-24</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>20.5,-34.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>19,-28</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>48.5,-22.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_INVERTER</type>
<position>33,-27.5</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>36.5,-32</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_OR2</type>
<position>55.5,-28</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>GA_LED</type>
<position>60.5,-28</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>46,-14</position>
<gparam>LABEL_TEXT 2x1 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>36.5,-37.5</position>
<gparam>LABEL_TEXT Using AOI logic</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-14,29.5,-14</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>29.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>29.5,-14,29.5,-14</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-14 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-17,27.5,-16</points>
<intersection>-17 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-16,29.5,-16</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-17,27.5,-17</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-12.5,31.5,-10.5</points>
<connection>
<GID>2</GID>
<name>SEL_0</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-10.5,31.5,-10.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-15,35.5,-15</points>
<connection>
<GID>10</GID>
<name>N_in0</name></connection>
<connection>
<GID>2</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21,-27.5,30,-27.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>21 4</intersection>
<intersection>25 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>21,-28,21,-27.5</points>
<intersection>-28 7</intersection>
<intersection>-27.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>25,-31,25,-27.5</points>
<intersection>-31 6</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>25,-31,33.5,-31</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>25 5</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>21,-28,21,-28</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>21 4</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-27.5,36,-23.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-23.5,45.5,-23.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-24,32.5,-21.5</points>
<intersection>-24 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-21.5,45.5,-21.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-24,32.5,-24</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-34.5,32,-33</points>
<intersection>-34.5 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-33,33.5,-33</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-34.5,32,-34.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-27,52,-22.5</points>
<intersection>-27 1</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-27,52.5,-27</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-22.5,52,-22.5</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-32,46,-29</points>
<intersection>-32 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-29,52.5,-29</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39.5,-32,46,-32</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-28,59.5,-28</points>
<connection>
<GID>26</GID>
<name>N_in0</name></connection>
<connection>
<GID>24</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>21.6705,6.8864,113.471,-38.4886</PageViewport>
<gate>
<ID>32</ID>
<type>AE_MUX_4x1</type>
<position>47,-16</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>13 </input>
<input>
<ID>IN_3</ID>12 </input>
<output>
<ID>OUT</ID>18 </output>
<input>
<ID>SEL_0</ID>17 </input>
<input>
<ID>SEL_1</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>35.5,-13</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>35.5,-15.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>35.5,-18</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>35.5,-20.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>42,-8</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>42,-5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>46</ID>
<type>GA_LED</type>
<position>52,-16</position>
<input>
<ID>N_in0</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>48,-23.5</position>
<gparam>LABEL_TEXT 4x1 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-13,44,-13</points>
<connection>
<GID>32</GID>
<name>IN_3</name></connection>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-15.5,40.5,-15</points>
<intersection>-15.5 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-15,44,-15</points>
<connection>
<GID>32</GID>
<name>IN_2</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-15.5,40.5,-15.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-18,40.5,-17</points>
<intersection>-18 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-17,44,-17</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-18,40.5,-18</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-20.5,40.5,-19</points>
<intersection>-20.5 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-19,44,-19</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-20.5,40.5,-20.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-11,47,-8</points>
<connection>
<GID>32</GID>
<name>SEL_1</name></connection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-8,47,-8</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-11,48,-5</points>
<connection>
<GID>32</GID>
<name>SEL_0</name></connection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-5,48,-5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-16,51,-16</points>
<connection>
<GID>46</GID>
<name>N_in0</name></connection>
<connection>
<GID>32</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>7.38751,-4.68125,99.1875,-50.0563</PageViewport>
<gate>
<ID>48</ID>
<type>BA_DECODER_2x4</type>
<position>40.5,-21.5</position>
<input>
<ID>ENABLE</ID>19 </input>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT_0</ID>25 </output>
<output>
<ID>OUT_1</ID>24 </output>
<output>
<ID>OUT_2</ID>23 </output>
<output>
<ID>OUT_3</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>32,-20</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_TOGGLE</type>
<position>32,-22.5</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_TOGGLE</type>
<position>32,-25</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>56</ID>
<type>GA_LED</type>
<position>47,-19.5</position>
<input>
<ID>N_in0</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>GA_LED</type>
<position>54.5,-21</position>
<input>
<ID>N_in0</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>GA_LED</type>
<position>53,-23.5</position>
<input>
<ID>N_in0</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>GA_LED</type>
<position>47,-28</position>
<input>
<ID>N_in0</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>38.5,-31</position>
<gparam>LABEL_TEXT 2x4 Decoder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-20,37.5,-20</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>37.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37.5,-20,37.5,-20</points>
<connection>
<GID>48</GID>
<name>ENABLE</name></connection>
<intersection>-20 1</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-22.5,35.5,-22</points>
<intersection>-22.5 2</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-22,37.5,-22</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-22.5,35.5,-22.5</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-25,35.5,-23</points>
<intersection>-25 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-23,37.5,-23</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-25,35.5,-25</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-20,44.5,-19.5</points>
<intersection>-20 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-19.5,46,-19.5</points>
<connection>
<GID>56</GID>
<name>N_in0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-20,44.5,-20</points>
<connection>
<GID>48</GID>
<name>OUT_3</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43.5,-21,53.5,-21</points>
<connection>
<GID>48</GID>
<name>OUT_2</name></connection>
<connection>
<GID>58</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-23.5,44.5,-22</points>
<intersection>-23.5 1</intersection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-23.5,52,-23.5</points>
<connection>
<GID>60</GID>
<name>N_in0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-22,44.5,-22</points>
<connection>
<GID>48</GID>
<name>OUT_1</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-28,43.5,-23</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-28,46,-28</points>
<connection>
<GID>64</GID>
<name>N_in0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>